module insert_sort #(
  )(
  );

endmodule
