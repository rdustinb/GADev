module selection_sort ();

endmodule
