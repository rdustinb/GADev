`define DLY_FOUR 7
`define MUX_FOUR_ONE 25
`define MUX_FOUR_TWO 73
`define MUX_FOUR_THREE 137
