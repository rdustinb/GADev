real2hex(3.141592653589793, working);
$display("The Hex fixed point value is: %08h", working);

