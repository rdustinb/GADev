`define DLY_ONE 13
`define RESET_ONE 8'h03
