`define DLY_THREE 9
`define RESET_THREE 8'h37
