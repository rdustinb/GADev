module shell_sort ();

endmodule
