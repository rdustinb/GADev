`define DLY_TWO 11
`define RESET_TWO 8'h15
